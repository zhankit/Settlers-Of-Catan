0
4 4 4 4 4 g c 
4 4 4 4 4 g c 
4 4 4 4 4 g c 
4 4 4 4 4 g c 
4 5 2 9 2 4 0 10 2 10 5 7 4 2 4 8 1 6 3 12 3 11 0 6 0 3 1 9 3 3 1 8 0 4 1 5 2 11 
